MACRO skullfet_inverter
  CLASS BLOCK ;
  FOREIGN skullfet_inverter ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.700 BY 14.300 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.800 6.700 14.300 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.000 6.700 0.500 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 12.700800 ;
    PORT
      LAYER met1 ;
        RECT 0.100 6.950 0.600 7.750 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.240000 ;
    PORT
      LAYER met1 ;
        RECT 6.100 6.950 6.600 7.750 ;
    END
  END A
  OBS
      LAYER pwell ;
        RECT 0.650 8.650 5.850 13.800 ;
      LAYER nwell ;
        RECT 0.650 0.500 5.850 6.200 ;
      LAYER li1 ;
        RECT 0.900 12.950 1.700 13.700 ;
        RECT 0.700 12.450 1.900 12.950 ;
        RECT 0.100 11.050 1.600 11.550 ;
        RECT 0.100 3.450 0.600 11.050 ;
        RECT 6.100 4.450 6.600 9.850 ;
        RECT 0.100 2.950 1.700 3.450 ;
        RECT 1.000 1.550 1.900 2.050 ;
        RECT 0.950 0.850 1.650 1.550 ;
      LAYER mcon ;
        RECT 0.800 12.600 1.050 12.850 ;
        RECT 0.200 7.000 0.500 7.800 ;
        RECT 6.200 7.000 6.500 7.800 ;
        RECT 1.050 1.650 1.300 1.850 ;
      LAYER met1 ;
        RECT 0.100 12.950 0.500 14.300 ;
        RECT 2.330 13.200 4.490 13.470 ;
        RECT 0.100 12.500 1.100 12.950 ;
        RECT 2.060 12.930 4.490 13.200 ;
        RECT 1.520 12.390 5.030 12.930 ;
        RECT 1.250 11.310 5.300 12.390 ;
        RECT 1.250 11.040 2.060 11.310 ;
        RECT 1.250 10.770 1.790 11.040 ;
        RECT 1.520 10.500 1.790 10.770 ;
        RECT 2.870 10.500 3.680 11.310 ;
        RECT 4.490 11.040 5.300 11.310 ;
        RECT 4.760 10.770 5.300 11.040 ;
        RECT 4.760 10.500 5.030 10.770 ;
        RECT 1.520 10.230 2.060 10.500 ;
        RECT 2.600 10.230 3.950 10.500 ;
        RECT 4.490 10.230 5.030 10.500 ;
        RECT 1.520 9.960 3.140 10.230 ;
        RECT 3.410 9.960 4.760 10.230 ;
        RECT 2.060 9.690 2.870 9.960 ;
        RECT 3.680 9.690 4.760 9.960 ;
        RECT 2.330 9.150 4.220 9.690 ;
        RECT 0.710 8.880 1.520 9.150 ;
        RECT 2.330 8.880 2.600 9.150 ;
        RECT 2.870 8.880 3.140 9.150 ;
        RECT 3.410 8.880 3.680 9.150 ;
        RECT 3.950 8.880 4.220 9.150 ;
        RECT 5.030 8.880 5.840 9.150 ;
        RECT 0.440 8.340 1.790 8.880 ;
        RECT 4.760 8.340 6.110 8.880 ;
        RECT 0.710 8.070 2.330 8.340 ;
        RECT 4.220 8.070 5.840 8.340 ;
        RECT 0.100 7.750 0.620 7.890 ;
        RECT 1.520 7.800 2.600 8.070 ;
        RECT 3.950 7.800 5.030 8.070 ;
        RECT 0.600 6.950 0.620 7.750 ;
        RECT 2.060 7.530 3.140 7.800 ;
        RECT 3.410 7.530 4.490 7.800 ;
        RECT 6.100 7.750 6.600 7.890 ;
        RECT 2.600 6.990 3.950 7.530 ;
        RECT 0.100 6.900 0.620 6.950 ;
        RECT 2.060 6.720 3.140 6.990 ;
        RECT 3.410 6.720 4.490 6.990 ;
        RECT 6.100 6.900 6.600 6.950 ;
        RECT 0.710 6.450 2.600 6.720 ;
        RECT 3.950 6.450 6.110 6.720 ;
        RECT 0.440 6.180 2.060 6.450 ;
        RECT 4.490 6.180 6.110 6.450 ;
        RECT 0.440 5.910 1.520 6.180 ;
        RECT 5.030 5.910 6.110 6.180 ;
        RECT 0.440 5.640 1.250 5.910 ;
        RECT 5.300 5.640 6.110 5.910 ;
        RECT 0.710 5.370 0.980 5.640 ;
        RECT 2.330 5.370 2.600 5.640 ;
        RECT 2.870 5.370 3.140 5.640 ;
        RECT 3.410 5.370 3.680 5.640 ;
        RECT 3.950 5.370 4.220 5.640 ;
        RECT 5.570 5.370 5.840 5.640 ;
        RECT 2.330 4.830 4.220 5.370 ;
        RECT 2.060 4.560 2.870 4.830 ;
        RECT 3.680 4.560 4.760 4.830 ;
        RECT 1.520 4.290 3.140 4.560 ;
        RECT 3.410 4.290 4.760 4.560 ;
        RECT 1.520 4.020 2.060 4.290 ;
        RECT 2.600 4.020 3.950 4.290 ;
        RECT 4.490 4.020 5.030 4.290 ;
        RECT 1.520 3.750 1.790 4.020 ;
        RECT 1.250 3.480 1.790 3.750 ;
        RECT 1.250 3.210 2.060 3.480 ;
        RECT 2.870 3.210 3.680 4.020 ;
        RECT 4.760 3.750 5.030 4.020 ;
        RECT 4.760 3.480 5.300 3.750 ;
        RECT 4.490 3.210 5.300 3.480 ;
        RECT 1.250 2.130 5.300 3.210 ;
        RECT 0.100 1.550 1.350 1.950 ;
        RECT 1.520 1.590 5.030 2.130 ;
        RECT 0.100 0.000 0.600 1.550 ;
        RECT 2.060 1.320 4.490 1.590 ;
        RECT 2.330 1.050 4.490 1.320 ;
      LAYER via ;
        RECT 0.150 13.850 0.450 14.250 ;
        RECT 0.150 0.050 0.550 0.450 ;
      LAYER met2 ;
        RECT 0.100 13.800 0.500 14.300 ;
        RECT 2.330 13.200 4.490 13.470 ;
        RECT 2.060 12.930 4.490 13.200 ;
        RECT 1.520 12.390 5.030 12.930 ;
        RECT 1.250 11.310 5.300 12.390 ;
        RECT 1.250 11.040 2.060 11.310 ;
        RECT 1.250 10.770 1.790 11.040 ;
        RECT 1.520 10.500 1.790 10.770 ;
        RECT 2.870 10.500 3.680 11.310 ;
        RECT 4.490 11.040 5.300 11.310 ;
        RECT 4.760 10.770 5.300 11.040 ;
        RECT 4.760 10.500 5.030 10.770 ;
        RECT 1.520 10.230 2.060 10.500 ;
        RECT 2.600 10.230 3.950 10.500 ;
        RECT 4.490 10.230 5.030 10.500 ;
        RECT 1.520 9.960 3.140 10.230 ;
        RECT 3.410 9.960 4.760 10.230 ;
        RECT 2.060 9.690 2.870 9.960 ;
        RECT 3.680 9.690 4.760 9.960 ;
        RECT 2.330 9.150 4.220 9.690 ;
        RECT 0.710 8.880 1.520 9.150 ;
        RECT 2.330 8.880 2.600 9.150 ;
        RECT 2.870 8.880 3.140 9.150 ;
        RECT 3.410 8.880 3.680 9.150 ;
        RECT 3.950 8.880 4.220 9.150 ;
        RECT 5.030 8.880 5.840 9.150 ;
        RECT 0.440 8.340 1.790 8.880 ;
        RECT 4.760 8.340 6.110 8.880 ;
        RECT 0.710 8.070 2.330 8.340 ;
        RECT 4.220 8.070 5.840 8.340 ;
        RECT 1.520 7.800 2.600 8.070 ;
        RECT 3.950 7.800 5.030 8.070 ;
        RECT 2.060 7.530 3.140 7.800 ;
        RECT 3.410 7.530 4.490 7.800 ;
        RECT 2.600 6.990 3.950 7.530 ;
        RECT 2.060 6.720 3.140 6.990 ;
        RECT 3.410 6.720 4.490 6.990 ;
        RECT 0.710 6.450 2.600 6.720 ;
        RECT 3.950 6.450 6.110 6.720 ;
        RECT 0.440 6.180 2.060 6.450 ;
        RECT 4.490 6.180 6.110 6.450 ;
        RECT 0.440 5.910 1.520 6.180 ;
        RECT 5.030 5.910 6.110 6.180 ;
        RECT 0.440 5.640 1.250 5.910 ;
        RECT 5.300 5.640 6.110 5.910 ;
        RECT 0.710 5.370 0.980 5.640 ;
        RECT 2.330 5.370 2.600 5.640 ;
        RECT 2.870 5.370 3.140 5.640 ;
        RECT 3.410 5.370 3.680 5.640 ;
        RECT 3.950 5.370 4.220 5.640 ;
        RECT 5.570 5.370 5.840 5.640 ;
        RECT 2.330 4.830 4.220 5.370 ;
        RECT 2.060 4.560 2.870 4.830 ;
        RECT 3.680 4.560 4.760 4.830 ;
        RECT 1.520 4.290 3.140 4.560 ;
        RECT 3.410 4.290 4.760 4.560 ;
        RECT 1.520 4.020 2.060 4.290 ;
        RECT 2.600 4.020 3.950 4.290 ;
        RECT 4.490 4.020 5.030 4.290 ;
        RECT 1.520 3.750 1.790 4.020 ;
        RECT 1.250 3.480 1.790 3.750 ;
        RECT 1.250 3.210 2.060 3.480 ;
        RECT 2.870 3.210 3.680 4.020 ;
        RECT 4.760 3.750 5.030 4.020 ;
        RECT 4.760 3.480 5.300 3.750 ;
        RECT 4.490 3.210 5.300 3.480 ;
        RECT 1.250 2.130 5.300 3.210 ;
        RECT 1.520 1.590 5.030 2.130 ;
        RECT 2.060 1.320 4.490 1.590 ;
        RECT 2.330 1.050 4.490 1.320 ;
        RECT 0.100 0.000 0.600 0.500 ;
      LAYER via2 ;
        RECT 0.150 13.850 0.450 14.250 ;
        RECT 0.150 0.050 0.550 0.450 ;
      LAYER met3 ;
        RECT 0.000 0.900 6.700 13.400 ;
  END
END skullfet_inverter
END LIBRARY

