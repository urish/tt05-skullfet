MACRO skullfet_nand
  CLASS BLOCK ;
  FOREIGN skullfet_nand ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.200 BY 14.310 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.374000 ;
    PORT
      LAYER met1 ;
        RECT 11.745 12.015 14.445 12.555 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.374000 ;
    PORT
      LAYER met1 ;
        RECT 1.755 2.835 4.455 3.375 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 17.714699 ;
    PORT
      LAYER met1 ;
        RECT 10.935 10.800 13.770 11.340 ;
    END
  END Y
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.000 16.200 0.400 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.700 16.200 1.100 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 10.935 6.345 16.200 10.125 ;
        RECT 5.670 5.265 16.200 6.345 ;
        RECT 5.670 1.080 10.530 5.265 ;
      LAYER li1 ;
        RECT 2.430 12.825 6.750 13.365 ;
        RECT 2.430 9.450 2.970 12.825 ;
        RECT 11.745 12.015 14.445 12.555 ;
        RECT 9.720 11.340 11.475 11.880 ;
        RECT 10.935 10.800 13.770 11.340 ;
        RECT 13.230 9.450 13.770 10.800 ;
        RECT 0.405 5.670 1.485 6.480 ;
        RECT 14.715 6.345 15.255 6.480 ;
        RECT 0.945 4.600 1.485 5.670 ;
        RECT 13.230 4.050 13.770 6.210 ;
        RECT 9.720 3.510 13.770 4.050 ;
        RECT 14.715 5.670 15.795 6.345 ;
        RECT 1.755 2.835 4.455 3.375 ;
        RECT 14.715 2.565 15.255 5.670 ;
        RECT 9.450 2.025 15.255 2.565 ;
        RECT 9.450 1.485 10.395 2.025 ;
      LAYER mcon ;
        RECT 11.820 12.090 12.210 12.480 ;
        RECT 13.980 12.090 14.370 12.480 ;
        RECT 11.010 10.875 11.400 11.265 ;
        RECT 13.305 10.875 13.695 11.265 ;
        RECT 1.000 4.700 1.400 5.100 ;
        RECT 1.830 2.910 2.220 3.300 ;
        RECT 3.990 2.910 4.380 3.300 ;
        RECT 11.745 2.025 12.150 2.565 ;
      LAYER met1 ;
        RECT 7.155 13.635 9.315 13.905 ;
        RECT 6.885 13.365 9.315 13.635 ;
        RECT 6.345 12.825 9.855 13.365 ;
        RECT 6.075 11.745 10.125 12.825 ;
        RECT 6.075 11.475 6.885 11.745 ;
        RECT 6.075 11.205 6.615 11.475 ;
        RECT 6.345 10.935 6.615 11.205 ;
        RECT 7.695 10.935 8.505 11.745 ;
        RECT 9.315 11.475 10.125 11.745 ;
        RECT 9.585 11.205 10.125 11.475 ;
        RECT 9.585 10.935 9.855 11.205 ;
        RECT 6.345 10.665 6.885 10.935 ;
        RECT 7.425 10.665 8.775 10.935 ;
        RECT 9.315 10.665 9.855 10.935 ;
        RECT 6.345 10.395 7.965 10.665 ;
        RECT 8.235 10.395 9.585 10.665 ;
        RECT 6.885 10.125 7.695 10.395 ;
        RECT 8.505 10.125 9.585 10.395 ;
        RECT 1.485 9.585 3.105 9.855 ;
        RECT 7.155 9.585 9.045 10.125 ;
        RECT 13.095 9.585 14.715 9.855 ;
        RECT 0.945 9.315 3.645 9.585 ;
        RECT 5.535 9.315 6.345 9.585 ;
        RECT 7.155 9.315 7.425 9.585 ;
        RECT 7.695 9.315 7.965 9.585 ;
        RECT 8.235 9.315 8.505 9.585 ;
        RECT 8.775 9.315 9.045 9.585 ;
        RECT 9.855 9.315 10.665 9.585 ;
        RECT 12.285 9.315 15.255 9.585 ;
        RECT 0.945 9.045 2.835 9.315 ;
        RECT 3.375 9.045 4.185 9.315 ;
        RECT 0.405 8.235 2.565 9.045 ;
        RECT 3.645 8.775 4.185 9.045 ;
        RECT 5.265 8.775 6.615 9.315 ;
        RECT 9.585 8.775 10.935 9.315 ;
        RECT 12.285 9.045 12.825 9.315 ;
        RECT 13.365 9.045 15.255 9.315 ;
        RECT 12.015 8.775 12.555 9.045 ;
        RECT 3.645 8.505 4.995 8.775 ;
        RECT 5.535 8.505 7.155 8.775 ;
        RECT 9.045 8.505 10.665 8.775 ;
        RECT 11.205 8.505 12.555 8.775 ;
        RECT 13.635 8.775 15.525 9.045 ;
        RECT 3.375 8.235 4.725 8.505 ;
        RECT 6.345 8.235 7.425 8.505 ;
        RECT 8.775 8.235 9.855 8.505 ;
        RECT 11.475 8.235 12.825 8.505 ;
        RECT 13.635 8.235 15.795 8.775 ;
        RECT 0.405 7.965 3.915 8.235 ;
        RECT 4.185 7.965 4.995 8.235 ;
        RECT 6.885 7.965 7.965 8.235 ;
        RECT 8.235 7.965 9.315 8.235 ;
        RECT 11.205 7.965 12.015 8.235 ;
        RECT 12.285 7.965 15.795 8.235 ;
        RECT 0.405 7.695 3.645 7.965 ;
        RECT 4.185 7.695 4.725 7.965 ;
        RECT 0.405 7.425 3.915 7.695 ;
        RECT 4.185 7.425 4.995 7.695 ;
        RECT 7.425 7.425 8.775 7.965 ;
        RECT 11.475 7.695 12.015 7.965 ;
        RECT 12.555 7.695 15.795 7.965 ;
        RECT 11.205 7.425 12.015 7.695 ;
        RECT 12.285 7.425 15.795 7.695 ;
        RECT 0.405 6.885 2.565 7.425 ;
        RECT 3.375 7.155 4.725 7.425 ;
        RECT 6.885 7.155 7.965 7.425 ;
        RECT 8.235 7.155 9.315 7.425 ;
        RECT 11.475 7.155 12.825 7.425 ;
        RECT 0.675 6.615 2.565 6.885 ;
        RECT 3.645 6.885 4.995 7.155 ;
        RECT 5.535 6.885 7.425 7.155 ;
        RECT 8.775 6.885 10.935 7.155 ;
        RECT 11.205 6.885 12.555 7.155 ;
        RECT 3.645 6.615 4.185 6.885 ;
        RECT 5.265 6.615 6.885 6.885 ;
        RECT 9.315 6.615 10.935 6.885 ;
        RECT 0.945 6.345 2.835 6.615 ;
        RECT 3.375 6.345 3.915 6.615 ;
        RECT 0.945 6.075 3.915 6.345 ;
        RECT 5.265 6.345 6.345 6.615 ;
        RECT 9.855 6.345 10.935 6.615 ;
        RECT 12.015 6.615 12.555 6.885 ;
        RECT 13.635 6.615 15.795 7.425 ;
        RECT 12.015 6.345 12.825 6.615 ;
        RECT 13.365 6.345 15.255 6.615 ;
        RECT 5.265 6.075 6.075 6.345 ;
        RECT 10.125 6.075 10.935 6.345 ;
        RECT 12.555 6.075 15.255 6.345 ;
        RECT 1.485 5.805 3.105 6.075 ;
        RECT 5.535 5.805 5.805 6.075 ;
        RECT 7.155 5.805 7.425 6.075 ;
        RECT 7.695 5.805 7.965 6.075 ;
        RECT 8.235 5.805 8.505 6.075 ;
        RECT 8.775 5.805 9.045 6.075 ;
        RECT 10.395 5.805 10.665 6.075 ;
        RECT 13.095 5.805 14.715 6.075 ;
        RECT 7.155 5.265 9.045 5.805 ;
        RECT 0.900 4.600 1.500 5.200 ;
        RECT 6.885 4.995 7.695 5.265 ;
        RECT 8.505 4.995 9.585 5.265 ;
        RECT 6.345 4.725 7.965 4.995 ;
        RECT 8.235 4.725 9.585 4.995 ;
        RECT 6.345 4.455 6.885 4.725 ;
        RECT 7.425 4.455 8.775 4.725 ;
        RECT 9.315 4.455 9.855 4.725 ;
        RECT 6.345 4.185 6.615 4.455 ;
        RECT 6.075 3.915 6.615 4.185 ;
        RECT 6.075 3.645 6.885 3.915 ;
        RECT 7.695 3.645 8.505 4.455 ;
        RECT 9.585 4.185 9.855 4.455 ;
        RECT 9.585 3.915 10.125 4.185 ;
        RECT 9.315 3.645 10.125 3.915 ;
        RECT 6.075 2.565 10.125 3.645 ;
        RECT 6.345 2.025 9.855 2.565 ;
        RECT 6.885 1.755 9.315 2.025 ;
        RECT 11.610 1.800 15.400 3.105 ;
        RECT 7.155 1.485 9.315 1.755 ;
      LAYER via ;
        RECT 0.950 4.650 1.450 5.150 ;
        RECT 14.750 2.050 15.250 2.550 ;
      LAYER met2 ;
        RECT 7.155 13.635 9.315 13.905 ;
        RECT 6.885 13.365 9.315 13.635 ;
        RECT 6.345 12.825 9.855 13.365 ;
        RECT 6.075 11.745 10.125 12.825 ;
        RECT 6.075 11.475 6.885 11.745 ;
        RECT 6.075 11.205 6.615 11.475 ;
        RECT 6.345 10.935 6.615 11.205 ;
        RECT 7.695 10.935 8.505 11.745 ;
        RECT 9.315 11.475 10.125 11.745 ;
        RECT 9.585 11.205 10.125 11.475 ;
        RECT 9.585 10.935 9.855 11.205 ;
        RECT 6.345 10.665 6.885 10.935 ;
        RECT 7.425 10.665 8.775 10.935 ;
        RECT 9.315 10.665 9.855 10.935 ;
        RECT 6.345 10.395 7.965 10.665 ;
        RECT 8.235 10.395 9.585 10.665 ;
        RECT 6.885 10.125 7.695 10.395 ;
        RECT 8.505 10.125 9.585 10.395 ;
        RECT 1.485 9.585 3.105 9.855 ;
        RECT 7.155 9.585 9.045 10.125 ;
        RECT 13.095 9.585 14.715 9.855 ;
        RECT 0.945 9.315 3.645 9.585 ;
        RECT 7.155 9.315 7.425 9.585 ;
        RECT 7.695 9.315 7.965 9.585 ;
        RECT 8.235 9.315 8.505 9.585 ;
        RECT 8.775 9.315 9.045 9.585 ;
        RECT 12.285 9.315 15.255 9.585 ;
        RECT 0.945 9.045 2.835 9.315 ;
        RECT 3.375 9.045 4.185 9.315 ;
        RECT 12.285 9.045 12.825 9.315 ;
        RECT 13.365 9.045 15.255 9.315 ;
        RECT 0.405 8.235 2.565 9.045 ;
        RECT 3.645 8.775 4.185 9.045 ;
        RECT 12.015 8.775 12.555 9.045 ;
        RECT 3.645 8.505 4.995 8.775 ;
        RECT 11.205 8.505 12.555 8.775 ;
        RECT 13.635 8.775 15.525 9.045 ;
        RECT 3.375 8.235 4.725 8.505 ;
        RECT 11.475 8.235 12.825 8.505 ;
        RECT 13.635 8.235 15.795 8.775 ;
        RECT 0.405 7.965 3.915 8.235 ;
        RECT 4.185 7.965 4.995 8.235 ;
        RECT 11.205 7.965 12.015 8.235 ;
        RECT 12.285 7.965 15.795 8.235 ;
        RECT 0.405 7.695 3.645 7.965 ;
        RECT 4.185 7.695 4.725 7.965 ;
        RECT 11.475 7.695 12.015 7.965 ;
        RECT 12.555 7.695 15.795 7.965 ;
        RECT 0.405 7.425 3.915 7.695 ;
        RECT 4.185 7.425 4.995 7.695 ;
        RECT 11.205 7.425 12.015 7.695 ;
        RECT 12.285 7.425 15.795 7.695 ;
        RECT 0.405 6.885 2.565 7.425 ;
        RECT 3.375 7.155 4.725 7.425 ;
        RECT 11.475 7.155 12.825 7.425 ;
        RECT 0.675 6.615 2.565 6.885 ;
        RECT 3.645 6.885 4.995 7.155 ;
        RECT 11.205 6.885 12.555 7.155 ;
        RECT 3.645 6.615 4.185 6.885 ;
        RECT 12.015 6.615 12.555 6.885 ;
        RECT 13.635 6.615 15.795 7.425 ;
        RECT 0.945 6.345 2.835 6.615 ;
        RECT 3.375 6.345 3.915 6.615 ;
        RECT 12.015 6.345 12.825 6.615 ;
        RECT 13.365 6.345 15.255 6.615 ;
        RECT 0.945 6.075 3.915 6.345 ;
        RECT 12.555 6.075 15.255 6.345 ;
        RECT 1.485 5.805 3.105 6.075 ;
        RECT 7.155 5.805 7.425 6.075 ;
        RECT 7.695 5.805 7.965 6.075 ;
        RECT 8.235 5.805 8.505 6.075 ;
        RECT 8.775 5.805 9.045 6.075 ;
        RECT 13.095 5.805 14.715 6.075 ;
        RECT 7.155 5.265 9.045 5.805 ;
        RECT 0.900 0.700 1.500 5.200 ;
        RECT 6.885 4.995 7.695 5.265 ;
        RECT 8.505 4.995 9.585 5.265 ;
        RECT 6.345 4.725 7.965 4.995 ;
        RECT 8.235 4.725 9.585 4.995 ;
        RECT 6.345 4.455 6.885 4.725 ;
        RECT 7.425 4.455 8.775 4.725 ;
        RECT 9.315 4.455 9.855 4.725 ;
        RECT 6.345 4.185 6.615 4.455 ;
        RECT 6.075 3.915 6.615 4.185 ;
        RECT 6.075 3.645 6.885 3.915 ;
        RECT 7.695 3.645 8.505 4.455 ;
        RECT 9.585 4.185 9.855 4.455 ;
        RECT 9.585 3.915 10.125 4.185 ;
        RECT 9.315 3.645 10.125 3.915 ;
        RECT 6.075 2.565 10.125 3.645 ;
        RECT 6.345 2.025 9.855 2.565 ;
        RECT 6.885 1.755 9.315 2.025 ;
        RECT 7.155 1.485 9.315 1.755 ;
        RECT 14.700 0.000 15.300 2.600 ;
      LAYER via2 ;
        RECT 0.950 0.750 1.450 1.050 ;
        RECT 14.750 0.050 15.250 0.350 ;
  END
END skullfet_nand
END LIBRARY

